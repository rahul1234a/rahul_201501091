`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ict_3rd_sem.
// Engineer: savriya rahul.
// Module Name:  inverse_matrix. 
// Project Name: inverse_matrix on fpga.
// rollno: 201501091.
//////////////////////////////////////////////////////////////////////////////////
module inverse_matrix(ran_acc_mem,start,clk,wr_st) ;
input start,clk;
output [31:0]ran_acc_mem;
output reg [31:0]wr_st;

wire flag;
wire swap_count,swap_flag;
wire [5:0]input_add_ram;
reg wr_stflag;
reg delay ;
reg [3:0]address_of_ram;
reg [31:0]output_ram,input_ram;
reg [31:0]temp_a;
reg [1:0] next_stage;
real a[0:4][0:9];
integer row = 0,column = 0;
real k;
reg rowtemp_a,columntemp_a;
reg r_add_flag;
reg s_fl;

initial
	begin
		next_stage = 2'b00;
		address_of_ram = 0;
		rowtemp_a = 0;
		r_add_flag = 0;
		s_fl = 1;
		wr_stflag = 0;
		delay = 0;
	end
	
random_acess_memory your_instance_name (
  .clka(clk), // input clka
  .wea(wr_stflag), // input [0 : 0] wea
  .addra(address_of_ram), // input [3 : 0] addra
  .dina(input_ram), // input [15 : 0] dina
  .douta(ran_acc_mem) // output [15 : 0] douta
);



always@(posedge clk)
	begin
		if(next_stage == 2'b00)
			if(delay == 0)
				begin
					delay = 1;
					address_of_ram = address_of_ram + 1'b1;
				end
			else
				begin
					temp_a = ran_acc_mem;
					a[row][column] =  ran_acc_mem;
	
			if(column < 10)
				begin
					if(column == 9)
						begin
						row = row + 1'b1;
						column = 0;
						end
				else
					column = column + 1;
				end
		if( row == 4)
		begin
			if(column == 9)
			begin
				next_stage = 2'b01;
			end
		end
		address_of_ram = address_of_ram + 1'b1;
	end
	else if(next_stage == 2'b01)
	begin
		
		if(a[0][0] != 32'b0)
		begin
			k = a[1][0] / a[0][0];
			wr_st = k;
			
			a[1][0] = a[1][0] - ((k)*a[0][0]);
			a[1][1] = a[1][1] - ((k)*a[0][1]);
			a[1][2] = a[1][2] - ((k)*a[0][2]);
			a[1][3] = a[1][3] - ((k)*a[0][3]);
			a[1][4] = a[1][4] - ((k)*a[0][4]);
			a[1][5] = a[1][5] - ((k)*a[0][5]);
			a[1][6] = a[1][6] - ((k)*a[0][6]);
			a[1][7] = a[1][7] - ((k)*a[0][7]);
			a[1][8] = a[1][8] - ((k)*a[0][8]);
			a[1][9] = a[1][9] - ((k)*a[0][9]);
		end
		if(a[0][0] != 0)
		begin
			k = a[2][0] / a[0][0];
			wr_st = k;
			a[1][0] = a[1][0] - ((k)*a[0][0]);
			a[1][1] = a[1][1] - ((k)*a[0][1]);
			a[1][2] = a[1][2] - ((k)*a[0][2]);
			a[1][3] = a[1][3] - ((k)*a[0][3]);
			a[1][4] = a[1][4] - ((k)*a[0][4]);
			a[1][5] = a[1][5] - ((k)*a[0][5]);
			a[1][6] = a[1][6] - ((k)*a[0][6]);
			a[1][7] = a[1][7] - ((k)*a[0][7]);
			a[1][8] = a[1][8] - ((k)*a[0][8]);
			a[1][9] = a[1][9] - ((k)*a[0][9]);
		end
		if(a[0][0] != 0)
		begin
		
			k = a[3][0] / a[0][0];
			a[1][0] = a[1][0] - ((k)*a[0][0]);
			a[1][1] = a[1][1] - ((k)*a[0][1]);
			a[1][2] = a[1][2] - ((k)*a[0][2]);
			a[1][3] = a[1][3] - ((k)*a[0][3]);
			a[1][4] = a[1][4] - ((k)*a[0][4]);
			a[1][5] = a[1][5] - ((k)*a[0][5]);
			a[1][6] = a[1][6] - ((k)*a[0][6]);
			a[1][7] = a[1][7] - ((k)*a[0][7]);
			a[1][8] = a[1][8] - ((k)*a[0][8]);
			a[1][9] = a[1][9] - ((k)*a[0][9]);
		end
		if(a[0][0] != 0)
		begin
			k = a[4][0] / a[0][0];
			wr_st = k;
			a[1][0] = a[1][0] - ((k)*a[0][0]);
			a[1][1] = a[1][1] - ((k)*a[0][1]);
			a[1][2] = a[1][2] - ((k)*a[0][2]);
			a[1][3] = a[1][3] - ((k)*a[0][3]);
			a[1][4] = a[1][4] - ((k)*a[0][4]);
			a[1][5] = a[1][5] - ((k)*a[0][5]);
			a[1][6] = a[1][6] - ((k)*a[0][6]);
			a[1][7] = a[1][7] - ((k)*a[0][7]);
			a[1][8] = a[1][8] - ((k)*a[0][8]);
			a[1][9] = a[1][9] - ((k)*a[0][9]);
		end
		if(a[1][1] != 0)
		begin
			k = a[2][1] / a[1][1];
			wr_st = k;
			a[2][0] = a[2][0] - ((k)*a[1][0]);
			a[2][1] = a[2][1] - ((k)*a[1][1]);
			a[2][2] = a[2][2] - ((k)*a[1][2]);
			a[2][3] = a[2][3] - ((k)*a[1][3]);
			a[2][4] = a[2][4] - ((k)*a[1][4]);
			a[2][5] = a[2][5] - ((k)*a[1][5]);
			a[2][6] = a[2][6] - ((k)*a[1][6]);
			a[2][7] = a[2][7] - ((k)*a[1][7]);
			a[2][8] = a[2][8] - ((k)*a[1][8]);
			a[2][9] = a[2][9] - ((k)*a[1][9]);
		end
		if(a[1][1] != 0)
		begin
			k = a[3][1] / a[1][1];
			wr_st = k;
			a[2][0] = a[2][0] - ((k)*a[1][0]);
			a[2][1] = a[2][1] - ((k)*a[1][1]);
			a[2][2] = a[2][2] - ((k)*a[1][2]);
			a[2][3] = a[2][3] - ((k)*a[1][3]);
			a[2][4] = a[2][4] - ((k)*a[1][4]);
			a[2][5] = a[2][5] - ((k)*a[1][5]);
			a[2][6] = a[2][6] - ((k)*a[1][6]);
			a[2][7] = a[2][7] - ((k)*a[1][7]);
			a[2][8] = a[2][8] - ((k)*a[1][8]);
			a[2][9] = a[2][9] - ((k)*a[1][9]);
		end
		if(a[1][1] != 0)
		begin
			k = a[4][1] / a[1][1];
			wr_st = k;
			a[2][0] = a[2][0] - ((k)*a[1][0]);
			a[2][1] = a[2][1] - ((k)*a[1][1]);
			a[2][2] = a[2][2] - ((k)*a[1][2]);
			a[2][3] = a[2][3] - ((k)*a[1][3]);
			a[2][4] = a[2][4] - ((k)*a[1][4]);
			a[2][5] = a[2][5] - ((k)*a[1][5]);
			a[2][6] = a[2][6] - ((k)*a[1][6]);
			a[2][7] = a[2][7] - ((k)*a[1][7]);
			a[2][8] = a[2][8] - ((k)*a[1][8]);
			a[2][9] = a[2][9] - ((k)*a[1][9]);
		end
		if(a[2][2] != 0)
		begin
			k = a[3][2] / a[2][2];
			wr_st = k;
			a[3][0] = a[3][0] - ((k)*a[2][0]);
			a[3][1] = a[3][1] - ((k)*a[2][1]);
			a[3][2] = a[3][2] - ((k)*a[2][2]);
			a[3][3] = a[3][3] - ((k)*a[2][3]);
			a[3][4] = a[3][4] - ((k)*a[2][4]);
			a[3][5] = a[3][5] - ((k)*a[2][5]);
			a[3][6] = a[3][6] - ((k)*a[2][6]);
			a[3][7] = a[3][7] - ((k)*a[2][7]);
			a[3][8] = a[3][8] - ((k)*a[2][8]);
			a[3][9] = a[3][9] - ((k)*a[2][9]);
		end
		if(a[2][2] != 0)
		begin
			k = a[4][2] / a[2][2];
			wr_st = k;
			a[3][0] = a[3][0] - ((k)*a[2][0]);
			a[3][1] = a[3][1] - ((k)*a[2][1]);
			a[3][2] = a[3][2] - ((k)*a[2][2]);
			a[3][3] = a[3][3] - ((k)*a[2][3]);
			a[3][4] = a[3][4] - ((k)*a[2][4]);
			a[3][5] = a[3][5] - ((k)*a[2][5]);
			a[3][6] = a[3][6] - ((k)*a[2][6]);
			a[3][7] = a[3][7] - ((k)*a[2][7]);
			a[3][8] = a[3][8] - ((k)*a[2][8]);
			a[3][9] = a[3][9] - ((k)*a[2][9]);
		end
		if(a[3][3] != 0)
		begin
			k = a[4][3] / a[3][3];
			wr_st = k;
			a[4][0] = a[4][0] - ((k)*a[3][0]);
			a[4][1] = a[4][1] - ((k)*a[3][1]);
			a[4][2] = a[4][2] - ((k)*a[3][2]);
			a[4][3] = a[4][3] - ((k)*a[3][3]);
			a[4][4] = a[4][4] - ((k)*a[3][4]);
			a[4][5] = a[4][5] - ((k)*a[3][5]);
			a[4][6] = a[4][6] - ((k)*a[3][6]);
			a[4][7] = a[4][7] - ((k)*a[3][7]);
			a[4][8] = a[4][8] - ((k)*a[3][8]);
			a[4][9] = a[4][9] - ((k)*a[3][9]);
		end
		next_stage = 2'b10;
		address_of_ram = 0;
		row = 3;
		column = 3;
	end
	else if(next_stage == 2'b10 )
	begin
	if(a[4][4] != 0)
		begin
			k = a[3][4] / a[4][4];
			wr_st = k;
			a[3][0] = a[3][0] - ((k)*a[4][0]);
			a[3][1] = a[3][1] - ((k)*a[4][1]);
			a[3][2] = a[3][2] - ((k)*a[4][2]);
			a[3][3] = a[3][3] - ((k)*a[4][3]);
			a[3][4] = a[3][4] - ((k)*a[4][4]);
			a[3][5] = a[3][5] - ((k)*a[4][5]);
			a[3][6] = a[3][6] - ((k)*a[4][6]);
			a[3][7] = a[3][7] - ((k)*a[4][7]);
			a[3][8] = a[3][8] - ((k)*a[4][8]);
		end
		if(a[4][4] != 0)
		begin
			k = a[2][4] / a[4][4];
			wr_st = k;
			a[2][0] = a[2][0] - ((k)*a[4][0]);
			a[2][1] = a[2][1] - ((k)*a[4][1]);
			a[2][2] = a[2][2] - ((k)*a[4][2]);
			a[2][3] = a[2][3] - ((k)*a[4][3]);
			a[2][4] = a[2][4] - ((k)*a[4][4]);
			a[2][5] = a[2][5] - ((k)*a[4][5]);
			a[2][6] = a[2][6] - ((k)*a[4][6]);
			a[2][7] = a[2][7] - ((k)*a[4][7]);
			a[2][8] = a[2][8] - ((k)*a[4][8]);
		end
		if(a[4][4] != 0)
		begin
			k = a[1][4] / a[4][4];
			wr_st = k;
			a[1][0] = a[1][0] - ((k)*a[4][0]);
			a[1][1] = a[1][1] - ((k)*a[4][1]);
			a[1][2] = a[1][2] - ((k)*a[4][2]);
			a[1][3] = a[1][3] - ((k)*a[4][3]);
			a[1][4] = a[1][4] - ((k)*a[4][4]);
			a[1][5] = a[1][5] - ((k)*a[4][5]);
			a[1][6] = a[1][6] - ((k)*a[4][6]);
			a[1][7] = a[1][7] - ((k)*a[4][7]);
			a[1][8] = a[1][8] - ((k)*a[4][8]);
		end
		if(a[4][4] != 0)
		begin
			k = a[0][4] / a[4][4];
			wr_st = k;
			a[0][0] = a[0][0] - ((k)*a[4][0]);
			a[0][1] = a[0][1] - ((k)*a[4][1]);
			a[0][2] = a[0][2] - ((k)*a[4][2]);
			a[0][3] = a[0][3] - ((k)*a[4][3]);
			a[0][4] = a[0][4] - ((k)*a[4][4]);
			a[0][5] = a[0][5] - ((k)*a[4][5]);
			a[0][6] = a[0][6] - ((k)*a[4][6]);
			a[0][7] = a[0][7] - ((k)*a[4][7]);
			a[0][8] = a[0][8] - ((k)*a[4][8]);
		end
		if(a[3][3] != 0)
		begin
			k = a[2][3] / a[3][3];
			wr_st = k;
			a[2][0] = a[2][0] - ((k)*a[3][0]);
			a[2][1] = a[2][1] - ((k)*a[3][1]);
			a[2][2] = a[2][2] - ((k)*a[3][2]);
			a[2][3] = a[2][3] - ((k)*a[3][3]);
			a[2][4] = a[2][4] - ((k)*a[3][4]);
			a[2][5] = a[2][5] - ((k)*a[3][5]);
			a[2][6] = a[2][6] - ((k)*a[3][6]);
			a[2][7] = a[2][7] - ((k)*a[3][7]);
			a[2][8] = a[2][8] - ((k)*a[3][8]);
		end
		if(a[3][3] != 0)
		begin
			k = a[1][3] / a[3][3];
			wr_st = k;
			a[1][0] = a[1][0] - ((k)*a[3][0]);
			a[1][1] = a[1][1] - ((k)*a[3][1]);
			a[1][2] = a[1][2] - ((k)*a[3][2]);
			a[1][3] = a[1][3] - ((k)*a[3][3]);
			a[1][4] = a[1][4] - ((k)*a[3][4]);
			a[1][5] = a[1][5] - ((k)*a[3][5]);
			a[1][6] = a[1][6] - ((k)*a[3][6]);
			a[1][7] = a[1][7] - ((k)*a[3][7]);
			a[1][8] = a[1][8] - ((k)*a[3][8]);
		end
		if(a[3][3] != 0)
		begin
			k = a[0][3] / a[3][3];
			wr_st = k;
			a[0][0] = a[0][0] - ((k)*a[3][0]);
			a[0][1] = a[0][1] - ((k)*a[3][1]);
			a[0][2] = a[0][2] - ((k)*a[3][2]);
			a[0][3] = a[0][3] - ((k)*a[3][3]);
			a[0][4] = a[0][4] - ((k)*a[3][4]);
			a[0][5] = a[0][5] - ((k)*a[3][5]);
			a[0][6] = a[0][6] - ((k)*a[3][6]);
			a[0][7] = a[0][7] - ((k)*a[3][7]);
			a[0][8] = a[0][8] - ((k)*a[3][8]);
		end
		if(a[2][2] != 0)
		begin
			k = a[1][2] / a[2][2];
			wr_st = k;
			a[1][0] = a[1][0] - ((k)*a[2][0]);
			a[1][1] = a[1][1] - ((k)*a[2][1]);
			a[1][2] = a[1][2] - ((k)*a[2][2]);
			a[1][3] = a[1][3] - ((k)*a[2][3]);
			a[1][4] = a[1][4] - ((k)*a[2][4]);
			a[1][5] = a[1][5] - ((k)*a[2][5]);
			a[1][6] = a[1][6] - ((k)*a[2][6]);
			a[1][7] = a[1][7] - ((k)*a[2][7]);
			a[1][8] = a[1][8] - ((k)*a[2][8]);
		end
		if(a[2][2] != 0)
		begin
			k = a[0][2] / a[2][2];
			wr_st = k;
			a[0][0] = a[0][0] - ((k)*a[2][0]);
			a[0][1] = a[0][1] - ((k)*a[2][1]);
			a[0][2] = a[0][2] - ((k)*a[2][2]);
			a[0][3] = a[0][3] - ((k)*a[2][3]);
			a[0][4] = a[0][4] - ((k)*a[2][4]);
			a[0][5] = a[0][5] - ((k)*a[2][5]);
			a[0][6] = a[0][6] - ((k)*a[2][6]);
			a[0][7] = a[0][7] - ((k)*a[2][7]);
			a[0][8] = a[0][8] - ((k)*a[2][8]);
		end
		if(a[1][1] != 0)
		begin
			k = a[0][1] / a[1][1];
			a[0][0] = a[0][0] - ((k)*a[1][0]);
			a[0][1] = a[0][1] - ((k)*a[1][1]);
			a[0][2] = a[0][2] - ((k)*a[1][2]);
			a[0][3] = a[0][3] - ((k)*a[1][3]);
			a[0][4] = a[0][4] - ((k)*a[1][4]);
			a[0][5] = a[0][5] - ((k)*a[1][5]);
			a[0][6] = a[0][6] - ((k)*a[1][6]);
			a[0][7] = a[0][7] - ((k)*a[1][7]);
			a[0][8] = a[0][8] - ((k)*a[1][8]);
		end
		address_of_ram = 0;
		wr_stflag = 1'b1;
		row = 0;
		column = 0;
		next_stage = 2'b11;
		input_ram =  a[row][column];
		row <= row + 1;
		column <= column + 1;
	end
	else if(next_stage == 2'b11 )
	begin
		input_ram =  a[row][column];
		wr_st = row;
		if(column < 10)
			begin
				if(column == 9)
				begin
					row = row + 1'b1;
					column = 0;
				end
				else
					column = column + 1;
			end
			if( row == 5)
			begin
				if(column == 0)
				begin
					$finish;
				end
			end
		address_of_ram = address_of_ram + 1;
	end
end




endmodule
